module helloworld;

initial begin
	$display("Hello world!");
end

endmodule